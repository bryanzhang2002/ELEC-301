CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 20 20 
10 13 13 10 20 13 20 20 14 20 
18 17 20 16 16 20 20 20 10 13 
20 18 11 
40 100 30 200 9
0 71 1920 864
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1920 864
9961490 0
0
6 Title:
5 Name:
0
0
0
17
7 Ground~
168 310 412 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8953 0 0
0
0
11 Signal Gen~
195 275 387 0 19 64
0 3 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 1028443341
20
1 1000 0 0.05 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
9 -50m/50mV
-32 -30 31 -22
2 V2
-7 -40 7 -32
0
0
38 %D %1 %2 DC 0 SIN(0 50m 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
4441 0 0
0
0
10 Capacitor~
219 371 363 0 2 5
0 4 5
0
0 0 336 0
4 10uF
-14 -18 14 -10
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3618 0 0
0
0
7 Ground~
168 396 413 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6153 0 0
0
0
7 Ground~
168 241 323 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5394 0 0
0
0
2 +V
167 428 414 0 1 3
0 6
0
0 0 54128 180
3 -5V
7 -2 28 6
3 VEE
7 -12 28 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7734 0 0
0
0
12 NPN Trans:B~
219 423 363 0 3 7
0 8 5 6
0
0 0 848 0
6 2N3904
9 4 51 12
2 Q3
19 -8 33 0
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
9914 0 0
0
0
7 Ground~
168 451 292 0 1 3
0 2
0
0 0 53360 90
0
4 GND1
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3747 0 0
0
0
2 +V
167 364 205 0 1 3
0 10
0
0 0 54128 0
2 5V
-8 -15 6 -7
3 VCC
-11 -25 10 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3549 0 0
0
0
12 NPN Trans:B~
219 301 294 0 3 7
0 12 9 8
0
0 0 848 0
6 2N3904
10 3 52 11
2 Q2
18 -11 32 -3
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
7931 0 0
0
0
12 NPN Trans:B~
219 437 293 0 3 7
0 11 2 8
0
0 0 848 512
6 2N3904
-53 3 -11 11
2 Q1
-40 -11 -26 -3
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
9325 0 0
0
0
11 Signal Gen~
195 193 299 0 19 64
0 7 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1203982336 0 1028443341
20
1 100000 0 0.05 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
9 -50m/50mV
-32 -30 31 -22
2 V1
-7 -40 7 -32
0
0
40 %D %1 %2 DC 0 SIN(0 50m 100k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
8903 0 0
0
0
9 Resistor~
219 335 363 0 2 5
0 3 4
0
0 0 368 0
2 2k
-7 -14 7 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3834 0 0
0
0
9 Resistor~
219 396 389 0 3 5
0 2 5 -1
0
0 0 368 90
4 200k
-32 -3 -4 5
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3363 0 0
0
0
9 Resistor~
219 428 243 0 4 5
0 11 10 0 1
0
0 0 880 90
2 1k
8 0 22 8
3 RC1
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7668 0 0
0
0
9 Resistor~
219 306 247 0 4 5
0 12 10 0 1
0
0 0 880 90
2 1k
8 0 22 8
3 RC2
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4718 0 0
0
0
9 Resistor~
219 253 294 0 2 5
0 7 9
0
0 0 880 0
2 50
-7 -14 7 -6
2 Rs
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3874 0 0
0
0
17
2 1 2 0 0 8192 0 2 1 0 0 3
306 392
310 392
310 406
1 1 3 0 0 8320 0 2 13 0 0 4
306 382
309 382
309 363
317 363
2 1 4 0 0 12416 0 13 3 0 0 4
353 363
347 363
347 363
362 363
2 0 5 0 0 4096 0 7 0 0 5 2
405 363
396 363
2 2 5 0 0 4224 0 3 14 0 0 3
380 363
396 363
396 371
1 1 2 0 0 0 0 4 14 0 0 2
396 407
396 407
1 3 6 0 0 4224 0 6 7 0 0 2
428 399
428 381
1 1 7 0 0 4224 0 12 17 0 0 2
224 294
235 294
2 1 2 0 0 4224 0 12 5 0 0 3
224 304
241 304
241 317
0 1 8 0 0 4096 0 0 7 12 0 2
428 319
428 345
1 2 2 0 0 0 0 8 11 0 0 2
444 293
451 293
3 3 8 0 0 8320 0 10 11 0 0 4
306 312
306 319
428 319
428 311
2 2 9 0 0 4224 0 17 10 0 0 2
271 294
283 294
2 0 10 0 0 8320 0 15 0 0 15 3
428 225
428 218
364 218
2 1 10 0 0 0 0 16 9 0 0 4
306 229
306 218
364 218
364 214
1 1 11 0 0 4224 0 15 11 0 0 2
428 261
428 275
1 1 12 0 0 4224 0 16 10 0 0 2
306 265
306 276
0
0
16 0 0
0
0
0
0 0 0
0
0 0 0
10 1 0.001 1e+011
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
2492404 8417856 100 100 0 0
77 66 1877 396
0 551 1920 1031
450 66
437 66
1877 284
1877 393
428 269
0.00103741 0.001 0.1 -3.88 0.005 0.005
12297 0
4 0.001 3
1
306 270
0 12 0 0 1	0 17 0 0
3146952 8550464 100 100 0 0
77 66 917 396
961 79 1921 559
917 66
77 66
917 66
917 396
0 0
4.94359e-315 0 4.94359e-315 0 4.94359e-315 4.94359e-315
12385 0
4 0.001 10
0
3934596 4618306 100 100 0 0
77 66 917 396
961 559 1921 1039
876 66
77 66
917 329
917 334
428 274
6.68125e-315 4.85009e-315 1.60899e-314 1.60958e-314 6.77444e-315 6.77444e-315
12435 0
4 3e+009 5e+009
1
266 131
0 10 0 0 1	0 17 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
