CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 20 20 
10 13 13 10 20 13 20 20 14 20 
18 17 20 16 16 20 20 20 10 13 
20 18 11 
610 150 30 200 9
1 79 961 1040
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
1 79 961 1040
9961490 0
0
6 Title:
5 Name:
0
0
0
16
11 Signal Gen~
195 968 511 0 64 64
0 3 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1203982336 0 981668463
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 -2118630188
20
1 100000 0 0.001 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
7 -1m/1mV
-25 -30 24 -22
2 V1
-5 -39 9 -31
0
0
39 %D %1 %2 DC 0 SIN(0 1m 100k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
8953 0 0
0
0
10 Capacitor~
219 771 374 0 2 5
0 7 2
0
0 0 848 90
7 0.027uF
3 6 52 14
2 CB
13 -7 27 1
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
4441 0 0
0
0
7 Ground~
168 905 505 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3618 0 0
0
0
2 +V
167 905 337 0 1 3
0 6
0
0 0 54128 0
3 12V
-10 -14 11 -6
3 VCC
-10 -25 11 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6153 0 0
0
0
12 NPN Trans:B~
219 900 425 0 3 7
0 6 8 4
0
0 0 848 0
6 2N3904
8 3 50 11
2 Q2
18 -9 32 -1
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
5394 0 0
0
0
12 NPN Trans:B~
219 737 418 0 3 7
0 8 7 5
0
0 0 848 270
6 2N3904
-22 18 20 26
2 Q1
-8 9 6 17
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
7734 0 0
0
0
10 Capacitor~
219 667 425 0 2 5
0 2 5
0
0 0 848 0
5 5.6uF
-18 -18 17 -10
3 CC1
-10 -28 11 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
9914 0 0
0
0
7 Ground~
168 670 366 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3747 0 0
0
0
10 Capacitor~
219 973 457 0 2 5
0 4 3
0
0 0 848 0
5 5.6uF
-16 -19 19 -11
3 CC2
-9 -29 12 -21
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3549 0 0
0
0
7 Ground~
168 646 453 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7931 0 0
0
0
7 Ground~
168 1006 541 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9325 0 0
0
0
9 Resistor~
219 735 379 0 4 5
0 7 2 0 -1
0
0 0 880 90
4 100k
3 2 31 10
3 RB2
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8903 0 0
0
0
9 Resistor~
219 829 378 0 4 5
0 7 6 0 1
0
0 0 880 90
4 150k
3 3 31 11
3 RB1
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3834 0 0
0
0
9 Resistor~
219 905 481 0 3 5
0 2 4 -1
0
0 0 880 90
4 6.8k
1 0 29 8
3 RE2
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3363 0 0
0
0
9 Resistor~
219 869 378 0 4 5
0 8 6 0 1
0
0 0 880 90
4 3.9k
3 2 31 10
3 RC1
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7668 0 0
0
0
9 Resistor~
219 694 382 0 4 5
0 5 2 0 -1
0
0 0 880 90
4 8.2k
5 0 33 8
3 RE1
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4718 0 0
0
0
19
2 1 2 0 0 8192 0 1 11 0 0 3
999 516
1006 516
1006 535
2 1 3 0 0 8336 0 9 1 0 0 4
982 457
1006 457
1006 506
999 506
1 1 2 0 0 8192 0 7 10 0 0 3
658 425
646 425
646 447
1 0 4 0 0 4224 0 9 0 0 5 2
964 457
905 457
3 2 4 0 0 0 0 5 14 0 0 2
905 443
905 463
2 0 2 0 0 8192 0 2 0 0 7 3
771 365
771 345
735 345
0 2 2 0 0 4224 0 0 12 8 0 3
683 345
735 345
735 361
1 2 2 0 0 0 0 8 16 0 0 4
670 360
670 345
694 345
694 364
2 0 5 0 0 4096 0 7 0 0 10 2
676 425
684 425
1 3 5 0 0 16512 0 16 6 0 0 5
694 400
694 425
684 425
684 425
717 425
2 0 6 0 0 8192 0 13 0 0 16 3
829 360
829 346
860 346
1 0 7 0 0 4096 0 2 0 0 13 2
771 383
771 403
1 1 7 0 0 8320 0 13 12 0 0 4
829 396
829 403
735 403
735 397
2 1 7 0 0 0 0 6 12 0 0 4
735 402
735 394
735 394
735 397
1 1 2 0 0 0 0 14 3 0 0 4
905 499
905 502
905 502
905 499
2 1 6 0 0 16384 0 15 4 0 0 5
869 360
869 346
860 346
860 346
905 346
1 0 8 0 0 4096 0 15 0 0 19 2
869 396
869 425
1 1 6 0 0 4224 0 5 4 0 0 2
905 407
905 346
1 2 8 0 0 4224 0 6 5 0 0 2
753 425
882 425
0
0
8 0 0
0
0
0
0 0 0
0
0 0 0
10 1 0.001 1e+013
0 5e-005 2e-007 2e-007
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
5243492 4356162 100 100 0 0
77 66 925 426
56 977 1026 1498
925 66
77 66
925 66
925 426
0 0
1e+013 0.001 0.3 -0.3 1e+013 1e+013
12435 0
5 3e+012 5e+012
1
1006 457
0 3 0 0 1	0 2 0 0
3148124 8550976 100 100 0 0
77 66 917 396
960 71 1920 551
917 66
77 66
917 66
917 396
0 0
5e-005 0 5e-005 0 5e-005 5e-005
12441 0
5 1e-005 10
0
6556012 4421696 100 100 0 0
77 66 917 396
960 551 1920 1031
917 66
77 66
917 66
917 66
0 0
4 1 0.0036 0 3 3
12401 0
4 1 2
1
581 461
0 5 0 0 2	0 20 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
