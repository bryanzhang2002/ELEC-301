CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 20 20 
10 13 13 10 20 13 20 20 14 20 
18 17 20 16 16 20 20 20 10 13 
20 18 11 
110 150 30 200 9
321 102 1268 965
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
321 102 1268 965
77070354 256
0
6 Title:
5 Name:
0
0
0
14
12 NPN Trans:B~
219 396 342 0 3 7
0 5 6 3
0
0 0 848 0
6 2N4401
18 0 60 8
2 Q1
32 -10 46 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
8953 0 0
0
0
7 Ground~
168 486 360 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4441 0 0
0
0
7 Ground~
168 369 414 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3618 0 0
0
0
10 Capacitor~
219 450 315 0 2 5
0 5 4
0
0 0 848 0
4 10uF
-14 -18 14 -10
3 CC2
-10 -28 11 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6153 0 0
0
0
10 Capacitor~
219 450 387 0 2 5
0 2 3
0
0 0 848 90
4 10uF
8 0 36 8
2 CE
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5394 0 0
0
0
2 +V
167 360 252 0 1 3
0 7
0
0 0 54128 0
3 15V
-9 -19 12 -11
3 VCC
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7734 0 0
0
0
10 Capacitor~
219 297 342 0 2 5
0 8 6
0
0 0 848 0
4 10uF
-14 -18 14 -10
3 CC1
-10 -28 11 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
9914 0 0
0
0
11 Signal Gen~
195 207 378 0 19 64
0 9 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1176256512 0 1008981771
20
1 10000 0 0.01 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
9 -10m/10mV
-32 -30 31 -22
2 V1
-7 -40 7 -32
0
0
39 %D %1 %2 DC 0 SIN(0 10m 10k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3747 0 0
0
0
9 Resistor~
219 486 333 0 3 5
0 2 4 -1
0
0 0 880 90
4 5.1k
5 3 33 11
2 RL
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3549 0 0
0
0
9 Resistor~
219 405 387 0 3 5
0 2 3 -1
0
0 0 880 90
4 4.3k
1 0 29 8
2 RE
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7931 0 0
0
0
9 Resistor~
219 405 288 0 4 5
0 5 7 0 1
0
0 0 880 90
4 5.1k
-34 2 -6 10
2 RC
-22 -10 -8 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9325 0 0
0
0
9 Resistor~
219 315 297 0 4 5
0 6 7 0 1
0
0 0 880 90
4 110k
3 0 31 8
3 RB1
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8903 0 0
0
0
9 Resistor~
219 315 378 0 3 5
0 2 6 -1
0
0 0 880 90
3 62k
5 0 26 8
3 RB2
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3834 0 0
0
0
9 Resistor~
219 261 342 0 2 5
0 9 8
0
0 0 880 0
2 50
-7 -14 7 -6
2 RS
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3363 0 0
0
0
17
2 0 2 0 0 8320 0 8 0 0 9 3
238 383
238 406
315 406
3 0 3 0 0 8192 0 1 0 0 7 3
401 360
401 362
405 362
1 1 2 0 0 0 0 2 9 0 0 4
486 354
486 357
486 357
486 351
2 2 4 0 0 4224 0 4 9 0 0 2
459 315
486 315
0 1 5 0 0 4224 0 0 4 11 0 2
405 315
441 315
0 1 2 0 0 0 0 0 5 8 0 3
405 406
450 406
450 396
2 2 3 0 0 8320 0 10 5 0 0 4
405 369
405 361
450 361
450 378
1 1 2 0 0 0 0 10 3 0 0 4
405 405
405 406
369 406
369 408
1 1 2 0 0 0 0 13 3 0 0 4
315 396
315 406
369 406
369 408
2 0 6 0 0 4224 0 1 0 0 14 2
378 342
315 342
1 1 5 0 0 0 0 11 1 0 0 5
405 306
405 305
405 305
405 324
401 324
1 2 7 0 0 8320 0 6 11 0 0 4
360 261
360 266
405 266
405 270
2 1 7 0 0 0 0 12 6 0 0 4
315 279
315 266
360 266
360 261
0 1 6 0 0 0 0 0 12 15 0 2
315 342
315 315
2 2 6 0 0 0 0 7 13 0 0 3
306 342
315 342
315 360
2 1 8 0 0 4224 0 14 7 0 0 2
279 342
288 342
1 1 9 0 0 4224 0 8 14 0 0 3
238 373
238 342
243 342
0
0
17 0 2
0
0
0
0 0 0
0
0 0 0
10 1 0.001 1e+011
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
7736124 1210432 100 100 0 0
0 0 0 0
13 76 174 146
0 66
0 66
1883 66
1883 876
0 0
0 0 0 0 0 0
12401 0
4 1 10
1
243 342
0 9 0 0 2	0 17 0 0
7341108 8812608 100 100 0 0
77 66 917 246
1 694 959 1031
917 66
77 66
917 69
917 246
0 0
0.005 0 10.7733 8.4 0.005 0.005
12401 0
4 0.001 10
1
406 315
0 5 0 0 1	0 5 0 0
0 0 100 100 0 0
77 66 1883 876
0 0 0 0
1883 66
77 66
1883 66
1883 876
0 0
1e+011 0.001 80 -141.778 1e+011 1e+011
12531 0
0 3e+010 5e+010
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
