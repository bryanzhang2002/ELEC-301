CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 20 20 
10 13 13 10 20 13 20 20 14 20 
18 17 20 16 16 20 20 20 10 13 
20 18 11 
100 170 30 200 9
1 79 961 1040
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
1 79 961 1040
9961491 0
0
6 Title:
5 Name:
0
0
0
13
7 Ground~
168 241 358 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8953 0 0
0
0
2 +V
167 368 418 0 1 3
0 4
0
0 0 54128 180
4 -15V
3 -2 31 6
3 VEE
7 -12 28 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4441 0 0
0
0
12 NPN Trans:B~
219 310 371 0 3 7
0 3 3 4
0
0 0 848 512
6 2N3904
-51 2 -9 10
2 Q4
-28 -9 -14 -1
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
3618 0 0
0
0
12 NPN Trans:B~
219 423 371 0 3 7
0 5 3 4
0
0 0 848 0
6 2N3904
9 4 51 12
2 Q3
19 -8 33 0
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
6153 0 0
0
0
7 Ground~
168 451 292 0 1 3
0 2
0
0 0 53360 90
0
4 GND1
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5394 0 0
0
0
2 +V
167 364 205 0 1 3
0 8
0
0 0 54128 0
3 15V
-11 -15 10 -7
3 VCC
-11 -25 10 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7734 0 0
0
0
12 NPN Trans:B~
219 301 294 0 3 7
0 10 7 5
0
0 0 848 0
6 2N3904
10 2 52 10
2 Q2
19 -13 33 -5
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
9914 0 0
0
0
12 NPN Trans:B~
219 437 293 0 3 7
0 9 2 5
0
0 0 848 512
6 2N3904
-53 3 -11 11
2 Q1
-40 -11 -26 -3
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
3747 0 0
0
0
11 Signal Gen~
195 202 299 0 19 64
0 6 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1203982336 0 1028443341
20
1 100000 0 0.05 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
9 -50m/50mV
-32 -30 31 -22
2 V1
-7 -40 7 -32
0
0
40 %D %1 %2 DC 0 SIN(0 50m 100k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3549 0 0
0
0
9 Resistor~
219 271 345 0 3 5
0 2 3 -1
0
0 0 880 0
4 6.8k
-14 -14 14 -6
4 Rref
-14 -24 14 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7931 0 0
0
0
9 Resistor~
219 428 243 0 4 5
0 9 8 0 1
0
0 0 880 90
3 10k
5 0 26 8
3 RC1
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9325 0 0
0
0
9 Resistor~
219 306 247 0 4 5
0 10 8 0 1
0
0 0 880 90
3 10k
5 0 26 8
3 RC2
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8903 0 0
0
0
9 Resistor~
219 261 294 0 2 5
0 6 7
0
0 0 880 0
2 50
-7 -14 7 -6
2 Rs
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3834 0 0
0
0
16
0 0 3 0 0 4096 0 0 0 4 8 3
301 345
333 345
333 371
2 0 2 0 0 8320 0 9 0 0 3 3
233 304
241 304
241 345
1 1 2 0 0 0 0 10 1 0 0 3
253 345
241 345
241 352
1 2 3 0 0 0 0 3 10 0 0 3
301 353
301 345
289 345
1 0 4 0 0 4096 0 2 0 0 6 3
368 403
368 397
367 397
3 3 4 0 0 8320 0 3 4 0 0 4
301 389
301 397
428 397
428 389
0 1 5 0 0 4096 0 0 4 10 0 2
428 319
428 353
2 2 3 0 0 4224 0 3 4 0 0 2
324 371
405 371
1 2 2 0 0 0 0 5 8 0 0 2
444 293
451 293
3 3 5 0 0 8320 0 7 8 0 0 4
306 312
306 319
428 319
428 311
1 1 6 0 0 12416 0 9 13 0 0 4
233 294
228 294
228 294
243 294
2 2 7 0 0 12416 0 13 7 0 0 4
279 294
276 294
276 294
283 294
2 0 8 0 0 8320 0 11 0 0 14 3
428 225
428 218
364 218
2 1 8 0 0 0 0 12 6 0 0 4
306 229
306 218
364 218
364 214
1 1 9 0 0 4224 0 11 8 0 0 2
428 261
428 275
1 1 10 0 0 4224 0 12 7 0 0 2
306 265
306 276
0
0
25 0 2
0
0
0
0 0 0
0
0 0 0
10 1 0.001 1e+011
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
2558708 1079360 100 100 0 0
77 66 1239 576
0 71 161 141
1239 66
77 66
1239 66
1239 576
428 274
1e+011 0.001 -100 -100 1e+011 300
12385 0
4 1 10
1
306 270
0 10 0 0 1	0 16 0 0
3146952 8550464 100 100 0 0
77 66 917 396
961 79 1921 559
917 66
77 66
917 66
917 396
0 0
0.005 0 0.005 0 0.005 0.005
12385 0
4 0.001 10
0
3934596 4618306 100 100 0 0
77 66 917 396
961 559 1921 1039
876 66
77 66
917 329
917 334
428 274
2.07332e+010 0.001 -39.0909 -43.6364 1e+011 1e+011
12435 0
4 3e+009 5e+009
1
306 271
0 10 0 0 1	0 16 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
