CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 20 20 
10 13 13 10 20 13 20 20 14 20 
18 17 20 16 16 20 20 20 10 13 
20 18 11 
60 290 30 200 9
0 71 960 1032
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 960 1032
1150812178 0
0
6 Title:
5 Name:
0
0
0
19
10 Capacitor~
219 419 494 0 2 5
0 2 3
0
0 0 33616 90
4 22uF
8 0 36 8
2 CE
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
8953 0 0
0
0
7 Ground~
168 454 401 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4441 0 0
0
0
10 Capacitor~
219 422 360 0 2 5
0 4 2
0
0 0 848 0
4 22uF
-14 -18 14 -10
3 CC2
-10 -28 11 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3618 0 0
0
0
7 Ground~
168 246 398 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6153 0 0
0
0
7 Ground~
168 197 508 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5394 0 0
0
0
10 Capacitor~
219 226 450 0 2 5
0 7 6
0
0 0 848 0
4 22uF
-14 -18 14 -10
3 CC1
-10 -28 11 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7734 0 0
0
0
11 Signal Gen~
195 166 479 0 19 64
0 7 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1176256512 0 1000593163
20
1 10000 0 0.005 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
7 -5m/5mV
-25 -30 24 -22
2 V1
-7 -40 7 -32
0
0
38 %D %1 %2 DC 0 SIN(0 5m 10k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
9914 0 0
0
0
10 Capacitor~
219 265 378 0 2 5
0 2 8
0
0 0 848 0
5 220uF
-18 -18 17 -10
2 CB
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3747 0 0
0
0
12 NPN Trans:B~
219 391 378 0 3 7
0 4 8 9
0
0 0 848 0
6 2N3904
10 4 52 12
2 Q2
21 -6 35 2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 1 0 0
1 Q
3549 0 0
0
0
12 NPN Trans:B~
219 391 450 0 3 7
0 9 5 3
0
0 0 848 0
6 2N3904
4 -4 46 4
2 Q1
16 -14 30 -6
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
7931 0 0
0
0
7 Ground~
168 342 520 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9325 0 0
0
0
2 +V
167 342 306 0 1 3
0 10
0
0 0 54128 0
3 20V
-10 -15 11 -7
3 VCC
-11 -27 10 -19
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8903 0 0
0
0
9 Resistor~
219 454 379 0 3 5
0 2 2 -1
0
0 0 880 90
3 50k
5 0 26 8
2 RL
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3834 0 0
0
0
9 Resistor~
219 269 450 0 2 5
0 6 5
0
0 0 880 0
4 3.3k
-14 -14 14 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3363 0 0
0
0
9 Resistor~
219 396 495 0 3 5
0 2 3 -1
0
0 0 880 90
4 2.4k
-33 0 -5 8
2 RE
-18 -12 -4 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7668 0 0
0
0
9 Resistor~
219 288 495 0 3 5
0 2 5 -1
0
0 0 880 90
3 51k
-25 0 -4 8
3 RB3
-25 -9 -4 -1
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4718 0 0
0
0
9 Resistor~
219 288 414 0 2 5
0 5 8
0
0 0 880 90
3 43k
5 1 26 9
3 RB2
6 -10 27 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3874 0 0
0
0
9 Resistor~
219 396 342 0 4 5
0 4 10 0 1
0
0 0 880 90
4 2.4k
-33 1 -5 9
2 RC
-20 -13 -6 -5
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6671 0 0
0
0
9 Resistor~
219 288 342 0 4 5
0 8 10 0 1
0
0 0 880 90
3 75k
5 4 26 12
3 RB1
4 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3789 0 0
0
0
23
2 1 2 0 0 8192 0 13 2 0 0 4
454 361
485 361
485 395
454 395
2 2 3 0 0 4224 0 15 1 0 0 3
396 477
419 477
419 485
1 1 2 0 0 0 0 1 15 0 0 3
419 503
419 513
396 513
1 1 2 0 0 0 0 2 13 0 0 4
454 395
454 398
454 398
454 397
2 2 2 0 0 128 0 3 13 0 0 3
431 360
454 360
454 361
1 1 4 0 0 4224 0 3 9 0 0 2
413 360
396 360
2 1 2 0 0 0 0 7 5 0 0 2
197 484
197 502
2 0 5 0 0 12288 0 14 0 0 17 4
287 450
284 450
284 450
288 450
2 1 6 0 0 4224 0 6 14 0 0 2
235 450
251 450
1 1 7 0 0 4240 0 7 6 0 0 3
197 474
197 450
217 450
1 1 2 0 0 0 0 8 4 0 0 3
256 378
246 378
246 392
0 2 8 0 0 4096 0 0 8 19 0 2
290 378
274 378
1 1 4 0 0 0 0 9 18 0 0 2
396 360
396 360
1 0 2 0 0 0 0 11 0 0 15 2
342 514
342 513
1 1 2 0 0 4224 0 16 15 0 0 2
288 513
396 513
3 2 3 0 0 0 0 10 15 0 0 2
396 468
396 477
2 0 5 0 0 4224 0 10 0 0 18 2
373 450
288 450
1 2 5 0 0 0 0 17 16 0 0 2
288 432
288 477
2 0 8 0 0 4224 0 9 0 0 20 2
373 378
288 378
1 2 8 0 0 0 0 19 17 0 0 2
288 360
288 396
3 1 9 0 0 4224 0 9 10 0 0 2
396 396
396 432
2 1 10 0 0 8320 0 19 12 0 0 3
288 324
288 315
342 315
1 2 10 0 0 0 0 12 18 0 0 3
342 315
396 315
396 324
0
0
25 0 2
0
0
0
0 0 0
0
0 0 0
10 1 0.001 1e+010
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
1902730 1210432 100 100 0 0
77 66 917 396
0 71 161 141
917 66
77 66
917 66
917 396
0 0
0.005 0 2.26381e-320 9.7224e-311 0.005 0.005
12401 0
4 1 10
1
396 326
0 10 0 0 2	18 0 0 0
2886116 8812608 100 100 0 0
77 66 917 396
960 71 1920 551
851 66
786 66
917 94
917 157
0 0
0.00460714 0.00422024 1.39636e-006 9.38182e-007 0.005 0.005
12409 0
4 0.001 10
1
219 450
0 7 0 0 1	6 0 0 0
4784876 4356672 100 100 0 0
77 66 922 396
960 551 1920 1031
922 66
77 66
922 229
922 333
0 0
1e+010 0.001 1.00364 0.816364 1e+010 1e+010
12435 0
4 3e+009 5e+009
1
203 450
0 7 0 0 2	0 10 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
