CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 20 20 
10 13 13 10 20 13 20 20 14 20 
18 17 20 16 16 20 20 20 10 13 
20 18 11 
200 140 30 200 9
30 99 990 1060
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
30 99 990 1060
77070354 256
0
6 Title:
5 Name:
0
0
0
15
7 Ground~
168 522 360 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8953 0 0
0
0
7 Ground~
168 513 441 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4441 0 0
0
0
7 Ground~
168 360 450 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3618 0 0
0
0
11 Signal Gen~
195 477 414 0 19 64
0 8 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 1050253722
20
1 1000 0 0.3 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
11 -300m/300mV
-40 31 37 39
2 V2
-6 22 8 30
0
0
39 %D %1 %2 DC 0 SIN(0 300m 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
6153 0 0
0
0
10 Capacitor~
219 441 369 0 2 5
0 5 9
0
0 0 848 0
4 10uF
-14 20 14 28
3 CC1
-10 11 11 19
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5394 0 0
0
0
10 Capacitor~
219 468 324 0 2 5
0 4 7
0
0 0 848 0
4 10uF
-14 -18 14 -10
3 CC2
-10 -28 11 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7734 0 0
0
0
2 +V
167 360 252 0 1 3
0 6
0
0 0 54128 0
3 15V
-9 -13 12 -5
3 VCC
-7 -24 14 -16
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
9914 0 0
0
0
12 NPN Trans:B~
219 396 351 0 3 7
0 4 3 5
0
0 0 848 0
7 2N2222A
8 0 57 8
2 Q1
9 -12 23 -4
0
0
14 %D %1 %2 %3 %M
0
0
5 TO-18
7

0 3 2 1 3 2 1 0
81 0 0 0 1 0 0 0
1 Q
3747 0 0
0
0
10 Capacitor~
219 279 387 0 2 5
0 2 3
0
0 0 848 90
4 10uF
-36 -1 -8 7
2 CB
-19 -11 -5 -3
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3549 0 0
0
0
9 Resistor~
219 486 369 0 2 5
0 9 8
0
0 0 880 0
2 50
-7 -14 7 -6
2 RS
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7931 0 0
0
0
9 Resistor~
219 522 342 0 3 5
0 2 7 -1
0
0 0 880 90
4 5.1k
3 0 31 8
2 R5
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9325 0 0
0
0
9 Resistor~
219 405 405 0 3 5
0 2 5 -1
0
0 0 880 90
4 4.3k
-27 -3 1 5
2 RE
-20 -15 -6 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8903 0 0
0
0
9 Resistor~
219 405 297 0 4 5
0 4 6 0 1
0
0 0 880 90
4 5.1k
4 1 32 9
2 RC
8 -9 22 -1
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3834 0 0
0
0
9 Resistor~
219 315 315 0 4 5
0 3 6 0 1
0
0 0 880 90
4 110k
6 2 34 10
3 RB1
7 -13 28 -5
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3363 0 0
0
0
9 Resistor~
219 315 387 0 3 5
0 2 3 -1
0
0 0 880 90
3 62k
5 0 26 8
3 RB2
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7668 0 0
0
0
18
1 0 3 0 0 4096 0 14 0 0 2 2
315 333
315 352
2 0 3 0 0 8192 0 9 0 0 6 3
279 378
279 352
315 352
1 0 2 0 0 4096 0 3 0 0 4 2
360 444
360 432
0 1 2 0 0 4240 0 0 12 12 0 3
314 432
405 432
405 423
1 0 4 0 0 4224 0 6 0 0 15 2
459 324
405 324
0 2 3 0 0 8320 0 0 8 9 0 3
315 352
315 351
378 351
0 1 5 0 0 8320 0 0 5 8 0 3
405 379
405 369
432 369
3 2 5 0 0 0 0 8 12 0 0 3
401 369
405 369
405 387
2 0 3 0 0 0 0 15 0 0 0 2
315 369
315 349
1 0 6 0 0 4096 0 7 0 0 11 2
360 261
360 270
2 2 6 0 0 8320 0 14 13 0 0 4
315 297
315 270
405 270
405 279
1 1 2 0 0 0 0 9 15 0 0 4
279 396
279 432
315 432
315 405
1 1 2 0 0 0 0 1 11 0 0 4
522 354
522 353
522 353
522 360
2 2 7 0 0 4224 0 6 11 0 0 2
477 324
522 324
1 1 4 0 0 0 0 8 13 0 0 3
401 333
405 333
405 315
2 1 2 0 0 0 0 4 2 0 0 3
508 419
513 419
513 435
2 1 8 0 0 8320 0 10 4 0 0 4
504 369
512 369
512 409
508 409
2 1 9 0 0 4224 0 5 10 0 0 2
450 369
468 369
0
0
25 0 2
0
0
0
0 0 0
0
0 0 0
10 1 0.001 1e+011
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
7211998 1079360 100 100 0 0
0 0 0 0
0 71 161 141
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12401 0
4 1 10
1
495 324
0 7 0 0 1	0 14 0 0
5442246 8550464 100 100 0 0
77 66 917 396
961 79 1921 559
917 66
77 66
917 66
917 396
0 0
0.005 0 0.005 0 0.005 0.005
12401 0
4 0.001 10
0
9243284 4325442 100 100 0 0
77 66 1883 876
-100 894 1820 1855
1883 66
77 66
1883 291
1883 790
0 0
1e+011 0.001 80 -141.778 1e+011 1e+011
12531 0
5 3e+010 5e+010
1
509 324
0 7 0 0 1	0 14 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
