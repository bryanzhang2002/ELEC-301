CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 20 20 
10 13 13 10 20 13 20 20 14 20 
18 17 20 16 16 20 20 20 10 13 
20 18 11 
150 280 30 260 9
0 71 1920 551
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1920 551
77070354 256
0
6 Title:
5 Name:
0
0
0
12
9 I Source~
198 450 333 0 2 5
0 2 6
0
0 0 17264 180
5 100mA
13 -1 48 7
2 Ib
23 -10 37 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
73 0 0 0 1 0 0 0
2 Is
8953 0 0
0
0
12 NPN Trans:B~
219 231 303 0 3 7
0 3 4 2
0
0 0 848 0
6 2N3904
18 0 60 8
2 Q3
32 -10 46 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
4441 0 0
0
0
9 V Source~
197 321 330 0 2 5
0 3 2
0
0 0 17008 0
2 5V
16 0 30 8
4 Vce2
10 -10 38 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
3618 0 0
0
0
7 Ground~
168 240 357 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6153 0 0
0
0
9 V Source~
197 168 330 0 2 5
0 4 2
0
0 0 17008 0
3 10V
13 0 34 8
4 Vbe2
10 -10 38 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
5394 0 0
0
0
12 NPN Trans:B~
219 509 306 0 3 7
0 5 6 2
0
0 0 848 0
6 2N3904
18 0 60 8
2 Q2
32 -10 46 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
7734 0 0
0
0
9 V Source~
197 599 333 0 2 5
0 5 2
0
0 0 17008 0
2 5V
16 0 30 8
4 Vce1
10 -10 38 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
9914 0 0
0
0
7 Ground~
168 518 360 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3747 0 0
0
0
9 V Source~
197 684 333 0 2 5
0 8 2
0
0 0 17008 0
3 10V
13 0 34 8
3 Vbe
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
3549 0 0
0
0
7 Ground~
168 756 360 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7931 0 0
0
0
9 V Source~
197 837 333 0 2 5
0 7 2
0
0 0 17008 0
2 5V
16 0 30 8
3 Vce
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
9325 0 0
0
0
12 NPN Trans:B~
219 747 306 0 3 7
0 7 8 2
0
0 0 848 0
6 2N3904
18 0 60 8
2 Q1
32 -10 46 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
8903 0 0
0
0
16
1 0 2 0 0 0 0 1 0 0 9 2
450 354
450 354
1 0 2 0 0 0 0 4 0 0 4 2
240 351
240 351
3 0 2 0 0 4096 0 2 0 0 4 2
236 321
236 351
2 2 2 0 0 4224 0 5 3 0 0 2
168 351
321 351
1 1 3 0 0 8320 0 3 2 0 0 3
321 309
321 285
236 285
1 2 4 0 0 8320 0 5 2 0 0 3
168 309
168 303
213 303
1 0 2 0 0 0 0 8 0 0 9 2
518 354
518 354
3 0 2 0 0 0 0 6 0 0 9 2
514 324
514 354
0 2 2 0 0 0 0 0 7 0 0 2
446 354
599 354
1 1 5 0 0 8320 0 7 6 0 0 3
599 312
599 288
514 288
2 2 6 0 0 8320 0 1 6 0 0 3
450 312
450 306
491 306
1 0 2 0 0 0 0 10 0 0 14 2
756 354
756 354
3 0 2 0 0 0 0 12 0 0 14 2
752 324
752 354
2 2 2 0 0 0 0 9 11 0 0 2
684 354
837 354
1 1 7 0 0 8320 0 11 12 0 0 3
837 312
837 288
752 288
1 2 8 0 0 8320 0 9 12 0 0 3
684 312
684 306
729 306
0
0
4 0 0
0
0
4 Vce2
0 6 0.02
4 Vbe2
0.55 0.7 0.01
3 0 1 4
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
4851970 2128448 100 100 0 0
77 66 1877 876
0 71 1920 1032
1877 66
77 66
1877 673
1877 876
0 0
6 0 0.00100741 -0.002 6 6
12441 0
5 1 5e+035
0
4982818 2259520 100 100 0 0
77 66 887 636
612 183 1559 917
751 66
212 66
887 228
887 240
0 0
5.3568e-315 5.26354e-315 4.96064e-315 4.95797e-315 5.36716e-315 5.36716e-315
12441 0
4 1 5e+035
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
