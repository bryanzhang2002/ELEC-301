CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
120 300 30 200 9
0 71 1920 663
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1920 663
9961490 0
0
6 Title:
5 Name:
0
0
0
11
2 +V
167 526 456 0 1 3
0 6
0
0 0 53616 692
3 15V
-12 1 9 9
2 V2
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8953 0 0
0
0
2 +V
167 526 402 0 1 3
0 7
0
0 0 53616 0
4 -15V
-13 -15 15 -7
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4441 0 0
0
0
7 Ground~
168 497 484 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3618 0 0
0
0
10 Capacitor~
219 430 418 0 2 5
0 5 8
0
0 0 848 0
5 0.5uF
-18 -18 17 -10
1 C
-4 -28 3 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6153 0 0
0
0
10 Capacitor~
219 374 418 0 2 5
0 4 5
0
0 0 848 0
5 0.5uF
-18 -18 17 -10
1 C
-4 -28 3 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5394 0 0
0
0
10 Capacitor~
219 321 418 0 2 5
0 3 4
0
0 0 848 0
5 0.5uF
-18 -18 17 -10
1 C
-4 -28 3 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7734 0 0
0
0
10 Op-Amp5:A~
219 526 424 0 5 11
0 2 9 6 7 3
0
0 0 848 692
5 UA741
12 4 47 12
2 U4
13 -14 27 -6
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 256 1 0 0 0
1 U
9914 0 0
0
0
9 Resistor~
219 524 366 0 2 5
0 3 9
0
0 0 880 180
5 14.6k
-17 -14 18 -6
3 R29
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3747 0 0
0
0
9 Resistor~
219 404 449 0 3 5
0 2 5 -1
0
0 0 880 90
3 500
5 0 26 8
1 R
11 -10 18 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3549 0 0
0
0
9 Resistor~
219 347 449 0 3 5
0 2 4 -1
0
0 0 880 90
3 500
5 0 26 8
1 R
11 -10 18 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7931 0 0
0
0
9 Resistor~
219 468 418 0 2 5
0 8 9
0
0 0 880 0
3 500
-10 -14 11 -6
1 R
-4 -24 3 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9325 0 0
0
0
14
1 1 3 0 0 12416 0 6 8 0 0 6
312 418
301 418
301 324
556 324
556 366
542 366
0 2 4 0 0 4096 0 0 6 8 0 2
347 418
330 418
1 0 2 0 0 4224 0 9 0 0 9 2
404 467
497 467
1 1 2 0 0 0 0 10 9 0 0 2
347 467
404 467
2 0 5 0 0 4096 0 9 0 0 6 2
404 431
404 418
2 1 5 0 0 4224 0 5 4 0 0 2
383 418
421 418
5 1 3 0 0 0 0 7 8 0 0 4
544 424
556 424
556 366
542 366
2 1 4 0 0 8320 0 10 5 0 0 3
347 431
347 418
365 418
1 1 2 0 0 0 0 7 3 0 0 3
508 430
497 430
497 478
1 3 6 0 0 4224 0 1 7 0 0 4
526 441
526 436
526 436
526 437
1 4 7 0 0 4224 0 2 7 0 0 4
526 411
526 408
526 408
526 411
2 1 8 0 0 12416 0 4 11 0 0 4
439 418
437 418
437 418
450 418
2 2 9 0 0 8320 0 8 7 0 0 4
506 366
500 366
500 418
508 418
2 2 9 0 0 0 0 11 7 0 0 2
486 418
508 418
0
0
16 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.1 5e-007 5e-007
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
4262092 8550976 100 100 0 0
77 66 1217 546
333 218 1595 863
123 66
167 66
1217 522
1217 306
0 0
0.00411324 0.00797662 0.00117559 0.00117564 0.1 0.1
12297 0
4 1e-006 10
1
556 419
0 3 0 0 2	0 7 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
