CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 180 30 200 9
1 79 1706 1040
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
1 79 1706 1040
1083703315 0
0
6 Title:
5 Name:
0
0
0
44
11 Signal Gen~
195 114 399 0 64 64
0 9 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 981668463
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 -1623938926
20
1 1000 0 0.001 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
7 -1m/1mV
-25 -30 24 -22
2 V2
-7 -40 7 -32
0
0
37 %D %1 %2 DC 0 SIN(0 1m 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
8953 0 0
0
0
7 Ground~
168 502 419 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4441 0 0
0
0
7 Ground~
168 341 449 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3618 0 0
0
0
2 +V
167 341 270 0 1 3
0 5
0
0 0 53616 0
3 15V
-10 -16 11 -8
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6153 0 0
0
0
10 Capacitor~
219 460 371 0 2 5
0 6 3
0
0 0 336 0
4 10uF
-14 -18 14 -10
2 C2
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5394 0 0
0
0
12 NPN Trans:B~
219 420 339 0 3 7
0 5 7 6
0
0 0 848 0
6 2N3904
18 0 60 8
2 Q2
32 -10 46 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
7734 0 0
0
0
12 NPN Trans:B~
219 336 366 0 3 7
0 7 8 2
0
0 0 848 0
6 2N3904
18 0 60 8
2 Q1
32 -10 46 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
9914 0 0
0
0
10 Capacitor~
219 229 366 0 2 5
0 4 8
0
0 0 336 0
4 10uF
-14 -18 14 -10
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3747 0 0
0
0
11 Signal Gen~
195 1100 388 0 64 64
0 16 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 981668463
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 -1623938926
20
1 1000 0 0.001 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
7 -1m/1mV
-25 -30 24 -22
2 V6
-7 -40 7 -32
0
0
37 %D %1 %2 DC 0 SIN(0 1m 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3549 0 0
0
0
7 Ground~
168 1488 408 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7931 0 0
0
0
7 Ground~
168 1327 438 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9325 0 0
0
0
2 +V
167 1327 259 0 1 3
0 12
0
0 0 53616 0
3 15V
-10 -16 11 -8
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8903 0 0
0
0
10 Capacitor~
219 1446 360 0 2 5
0 13 10
0
0 0 336 0
4 10uF
-14 -18 14 -10
2 C6
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3834 0 0
0
0
12 NPN Trans:B~
219 1406 328 0 3 7
0 12 14 13
0
0 0 848 0
6 2N3904
18 0 60 8
2 Q6
32 -10 46 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
3363 0 0
0
0
12 NPN Trans:B~
219 1322 355 0 3 7
0 14 15 2
0
0 0 848 0
6 2N3904
18 0 60 8
2 Q5
32 -10 46 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
7668 0 0
0
0
10 Capacitor~
219 1215 355 0 2 5
0 11 15
0
0 0 336 0
4 10uF
-14 -18 14 -10
2 C5
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
4718 0 0
0
0
10 Capacitor~
219 740 358 0 2 5
0 18 22
0
0 0 336 0
4 10uF
-14 -18 14 -10
2 C4
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3874 0 0
0
0
12 NPN Trans:B~
219 847 358 0 3 7
0 21 22 2
0
0 0 848 0
6 2N3904
18 0 60 8
2 Q4
32 -10 46 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
6671 0 0
0
0
12 NPN Trans:B~
219 931 331 0 3 7
0 19 21 20
0
0 0 848 0
6 2N3904
18 0 60 8
2 Q3
32 -10 46 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
3789 0 0
0
0
10 Capacitor~
219 971 363 0 2 5
0 20 17
0
0 0 336 0
4 10uF
-14 -18 14 -10
2 C3
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
4871 0 0
0
0
2 +V
167 852 262 0 1 3
0 19
0
0 0 53616 0
3 15V
-10 -16 11 -8
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3750 0 0
0
0
7 Ground~
168 852 441 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8778 0 0
0
0
7 Ground~
168 1013 411 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
538 0 0
0
0
11 Signal Gen~
195 625 391 0 64 64
0 23 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 981668463
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 -1623938926
20
1 1000 0 0.001 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
7 -1m/1mV
-25 -30 24 -22
2 V3
-7 -40 7 -32
0
0
37 %D %1 %2 DC 0 SIN(0 1m 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
6843 0 0
0
0
9 Resistor~
219 502 398 0 3 5
0 2 3 -1
0
0 0 880 90
3 10k
5 0 26 8
3 RL3
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3136 0 0
0
0
9 Resistor~
219 425 398 0 3 5
0 2 6 -1
0
0 0 368 90
3 560
5 0 26 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5950 0 0
0
0
9 Resistor~
219 341 308 0 4 5
0 7 5 0 1
0
0 0 880 90
5 10.1k
4 0 39 8
3 RC3
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5670 0 0
0
0
9 Resistor~
219 267 320 0 4 5
0 8 5 0 1
0
0 0 368 90
4 330k
6 -4 34 4
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6828 0 0
0
0
9 Resistor~
219 267 398 0 3 5
0 2 8 -1
0
0 0 880 90
3 20k
5 0 26 8
3 RB2
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6735 0 0
0
0
9 Resistor~
219 171 366 0 2 5
0 4 9
0
0 0 368 180
2 5k
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8365 0 0
0
0
9 Resistor~
219 1358 465 0 2 5
0 11 10
0
0 0 880 0
5 10Meg
-18 -14 17 -6
3 Rf2
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4132 0 0
0
0
9 Resistor~
219 1488 387 0 3 5
0 2 10 -1
0
0 0 880 90
3 10k
5 0 26 8
3 RL2
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4551 0 0
0
0
9 Resistor~
219 1411 387 0 3 5
0 2 13 -1
0
0 0 368 90
3 560
5 0 26 8
2 R9
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3635 0 0
0
0
9 Resistor~
219 1327 297 0 4 5
0 14 12 0 1
0
0 0 880 90
3 10k
5 0 26 8
3 RC2
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3973 0 0
0
0
9 Resistor~
219 1253 309 0 4 5
0 15 12 0 1
0
0 0 368 90
4 330k
6 -4 34 4
2 R8
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3851 0 0
0
0
9 Resistor~
219 1253 387 0 3 5
0 2 15 -1
0
0 0 880 90
3 20k
5 0 26 8
3 RB3
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8383 0 0
0
0
9 Resistor~
219 1157 355 0 2 5
0 11 16
0
0 0 368 180
2 5k
-7 -14 7 -6
2 R7
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9334 0 0
0
0
9 Resistor~
219 682 358 0 2 5
0 18 23
0
0 0 368 180
2 5k
-7 -14 7 -6
2 R6
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7471 0 0
0
0
9 Resistor~
219 778 390 0 3 5
0 2 22 -1
0
0 0 880 90
3 20k
5 0 26 8
3 RB1
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3334 0 0
0
0
9 Resistor~
219 778 312 0 4 5
0 22 19 0 1
0
0 0 368 90
4 330k
6 -4 34 4
2 R5
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3559 0 0
0
0
9 Resistor~
219 852 300 0 4 5
0 21 19 0 1
0
0 0 880 90
3 10k
5 0 26 8
3 RC1
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
984 0 0
0
0
9 Resistor~
219 936 390 0 3 5
0 2 20 -1
0
0 0 368 90
3 560
5 0 26 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7557 0 0
0
0
9 Resistor~
219 1013 390 0 3 5
0 2 17 -1
0
0 0 880 90
3 10k
5 0 26 8
3 RL1
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3146 0 0
0
0
9 Resistor~
219 883 468 0 2 5
0 18 17
0
0 0 880 0
4 1Meg
-14 -14 14 -6
3 Rf1
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5687 0 0
0
0
60
0 0 3 0 0 8320 0 0 0 0 5 3
391 476
476 476
476 371
0 0 4 0 0 4224 0 0 0 0 19 3
355 476
202 476
202 366
0 1 5 0 0 4224 0 0 6 16 0 3
340 280
425 280
425 321
1 1 2 0 0 4096 0 2 25 0 0 4
502 413
502 419
502 419
502 416
2 2 3 0 0 0 0 5 25 0 0 3
469 371
502 371
502 380
1 0 6 0 0 4224 0 5 0 0 8 2
451 371
425 371
1 1 2 0 0 8192 0 3 26 0 0 4
341 443
341 435
425 435
425 416
3 2 6 0 0 0 0 6 26 0 0 2
425 357
425 380
2 0 7 0 0 4224 0 6 0 0 15 2
402 339
341 339
1 0 2 0 0 0 0 29 0 0 11 2
267 416
267 435
2 1 2 0 0 8320 0 1 3 0 0 4
145 404
145 435
341 435
341 443
3 1 2 0 0 0 0 7 3 0 0 2
341 384
341 443
2 0 8 0 0 4096 0 29 0 0 14 2
267 380
267 366
1 0 8 0 0 4096 0 28 0 0 18 2
267 338
267 366
1 1 7 0 0 0 0 27 7 0 0 2
341 326
341 348
1 2 5 0 0 0 0 4 27 0 0 6
341 279
341 280
340 280
340 280
341 280
341 290
2 1 5 0 0 0 0 28 4 0 0 4
267 302
267 280
341 280
341 279
2 2 8 0 0 4224 0 8 7 0 0 2
238 366
318 366
1 1 4 0 0 0 0 30 8 0 0 2
189 366
220 366
1 2 9 0 0 4224 0 1 30 0 0 3
145 394
145 366
153 366
2 0 10 0 0 8320 0 31 0 0 25 3
1376 465
1462 465
1462 360
1 0 11 0 0 4224 0 31 0 0 39 3
1340 465
1188 465
1188 355
0 1 12 0 0 4224 0 0 14 36 0 3
1326 269
1411 269
1411 310
1 1 2 0 0 0 0 10 32 0 0 4
1488 402
1488 408
1488 408
1488 405
2 2 10 0 0 0 0 13 32 0 0 3
1455 360
1488 360
1488 369
1 0 13 0 0 4224 0 13 0 0 28 2
1437 360
1411 360
1 1 2 0 0 0 0 11 33 0 0 4
1327 432
1327 424
1411 424
1411 405
3 2 13 0 0 0 0 14 33 0 0 2
1411 346
1411 369
2 0 14 0 0 4224 0 14 0 0 35 2
1388 328
1327 328
1 0 2 0 0 0 0 36 0 0 31 2
1253 405
1253 424
2 1 2 0 0 0 0 9 11 0 0 4
1131 393
1131 424
1327 424
1327 432
3 1 2 0 0 0 0 15 11 0 0 2
1327 373
1327 432
2 0 15 0 0 4096 0 36 0 0 34 2
1253 369
1253 355
1 0 15 0 0 4096 0 35 0 0 38 2
1253 327
1253 355
1 1 14 0 0 0 0 34 15 0 0 2
1327 315
1327 337
1 2 12 0 0 0 0 12 34 0 0 6
1327 268
1327 269
1326 269
1326 269
1327 269
1327 279
2 1 12 0 0 0 0 35 12 0 0 4
1253 291
1253 269
1327 269
1327 268
2 2 15 0 0 4224 0 16 15 0 0 2
1224 355
1304 355
1 1 11 0 0 0 0 37 16 0 0 2
1175 355
1206 355
1 2 16 0 0 4224 0 9 37 0 0 3
1131 383
1131 355
1139 355
2 0 17 0 0 8320 0 44 0 0 45 3
901 468
987 468
987 363
1 0 18 0 0 4224 0 44 0 0 59 3
865 468
713 468
713 358
0 1 19 0 0 4224 0 0 19 56 0 3
851 272
936 272
936 313
1 1 2 0 0 0 0 23 43 0 0 4
1013 405
1013 411
1013 411
1013 408
2 2 17 0 0 0 0 20 43 0 0 3
980 363
1013 363
1013 372
1 0 20 0 0 4224 0 20 0 0 48 2
962 363
936 363
1 1 2 0 0 0 0 22 42 0 0 4
852 435
852 427
936 427
936 408
3 2 20 0 0 0 0 19 42 0 0 2
936 349
936 372
2 0 21 0 0 4224 0 19 0 0 55 2
913 331
852 331
1 0 2 0 0 0 0 39 0 0 51 2
778 408
778 427
2 1 2 0 0 0 0 24 22 0 0 4
656 396
656 427
852 427
852 435
3 1 2 0 0 0 0 18 22 0 0 2
852 376
852 435
2 0 22 0 0 4096 0 39 0 0 54 2
778 372
778 358
1 0 22 0 0 4096 0 40 0 0 58 2
778 330
778 358
1 1 21 0 0 0 0 41 18 0 0 2
852 318
852 340
1 2 19 0 0 0 0 21 41 0 0 6
852 271
852 272
851 272
851 272
852 272
852 282
2 1 19 0 0 0 0 40 21 0 0 4
778 294
778 272
852 272
852 271
2 2 22 0 0 4224 0 17 18 0 0 2
749 358
829 358
1 1 18 0 0 0 0 38 17 0 0 2
700 358
731 358
1 2 23 0 0 4224 0 24 38 0 0 3
656 386
656 358
664 358
0
0
25 0 2
0
0
0
0 0 0
0
0 0 0
10 1 0.01 1e+008
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
722474 1079360 100 100 0 0
0 0 0 0
0 71 161 141
0 66
0 66
1217 66
1217 546
0 0
0 0 0 0 0 0
12401 0
4 1 10
1
491 371
0 3 0 0 1	0 5 0 0
1902902 8550464 100 100 0 0
77 66 917 396
696 693 1656 1173
917 66
77 66
917 66
917 396
0 0
0.005 0 0.005 0 0.005 0.005
12385 0
4 0.001 10
0
723260 4421696 978 1157 770 645
77 66 1887 876
0 71 1920 1032
1652 66
1652 66
1887 160
1887 361
0 0
1392.02 1392.02 44.7236 42.1499 1e+008 1e+008
45075 0
4 0.03 5
1
493 371
0 3 0 0 1	0 5 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
