CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 20 20 
10 13 13 10 20 13 20 20 14 20 
18 17 20 16 16 20 20 20 10 13 
20 18 11 
370 270 30 200 9
0 71 1920 1032
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1920 1032
211288082 256
0
6 Title:
5 Name:
0
0
0
17
12 V->I Source~
200 781 346 0 4 9
0 3 2 5 2
0
0 0 17232 0
3 0.1
-10 -12 11 -4
3 GV1
39 -3 60 5
0
0
17 %D %1 %2 %3 %4 %V
0
0
0
9

0 3 4 1 2 3 4 1 2 0
71 0 0 0 1 0 0 0
4 VcIs
8953 0 0
0
0
7 Ground~
168 655 382 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4441 0 0
0
0
7 Ground~
168 700 382 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3618 0 0
0
0
7 Ground~
168 763 382 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6153 0 0
0
0
7 Ground~
168 799 382 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5394 0 0
0
0
7 Ground~
168 853 382 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7734 0 0
0
0
7 Ground~
168 898 382 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9914 0 0
0
0
7 Ground~
168 565 382 0 1 3
0 2
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3747 0 0
0
0
10 Capacitor~
219 637 310 0 2 5
0 6 5
0
0 0 848 0
3 1uF
-11 -18 10 -10
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3549 0 0
0
0
11 Signal Gen~
195 529 346 0 64 64
0 7 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 1065353216
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 150867206
20
1 1000 0 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
5 -1/1V
-18 -30 17 -22
2 V2
-7 -40 7 -32
0
0
36 %D %1 %2 DC 0 SIN(0 1 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
7931 0 0
0
0
10 Capacitor~
219 700 346 0 2 5
0 2 5
0
0 0 848 90
4 10pF
8 0 36 8
2 C2
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
9325 0 0
0
0
10 Capacitor~
219 781 310 0 2 5
0 5 3
0
0 0 848 0
3 2pF
-11 -18 10 -10
2 C3
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
8903 0 0
0
0
10 Capacitor~
219 871 310 0 2 5
0 3 4
0
0 0 848 0
3 1uF
-11 -18 10 -10
2 C4
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3834 0 0
0
0
9 Resistor~
219 592 310 0 2 5
0 7 6
0
0 0 880 0
2 50
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3363 0 0
0
0
9 Resistor~
219 655 346 0 3 5
0 2 5 -1
0
0 0 880 90
2 1k
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7668 0 0
0
0
9 Resistor~
219 853 346 0 3 5
0 2 3 -1
0
0 0 880 90
2 4k
8 0 22 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4718 0 0
0
0
9 Resistor~
219 898 346 0 3 5
0 2 8 -1
0
0 0 880 90
2 4k
8 0 22 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3874 0 0
0
0
18
1 0 3 0 0 4112 0 1 0 0 4 2
801 319
801 310
2 0 3 0 0 4112 0 16 0 0 4 2
853 328
853 310
2 0 4 0 0 4240 0 13 0 0 0 2
880 310
898 310
2 1 3 0 0 4240 0 12 13 0 0 2
790 310
862 310
1 1 2 0 0 4112 0 3 11 0 0 2
700 376
700 355
3 0 5 0 0 4112 0 1 0 0 9 2
761 319
761 310
2 0 5 0 0 4112 0 11 0 0 9 2
700 337
700 310
2 0 5 0 0 16 0 15 0 0 9 2
655 328
655 310
2 1 5 0 0 4240 0 9 12 0 0 2
646 310
772 310
2 1 6 0 0 4240 0 14 9 0 0 2
610 310
628 310
2 1 2 0 0 8336 0 10 8 0 0 3
560 351
565 351
565 376
1 1 7 0 0 4240 0 10 14 0 0 3
560 341
560 310
574 310
4 1 2 0 0 16 0 1 4 0 0 3
761 373
761 376
763 376
1 1 2 0 0 16 0 7 17 0 0 4
898 376
898 361
898 361
898 364
2 1 2 0 0 16 0 1 5 0 0 3
801 373
801 376
799 376
1 1 2 0 0 16 0 6 16 0 0 4
853 376
853 361
853 361
853 364
1 1 2 0 0 16 0 2 15 0 0 4
655 376
655 361
655 361
655 364
2 0 8 0 0 4240 0 17 0 0 0 2
898 328
898 310
0
0
8 0 0
0
0
0
0 0 0
0
0 0 0
10 1 0.01 1e+011
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
1116612 4421696 100 100 0 0
77 66 1884 576
5 370 1925 1023
1884 66
77 66
1884 67
1884 516
0 0
1e+011 0.01 -0.470588 -211.294 1e+011 1e+011
12435 0
5 3e+010 5e+010
1
529 346
0 0 0 0 0	10 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
