CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 20 20 
10 13 13 10 20 13 20 20 14 20 
18 17 20 16 16 20 20 20 10 13 
20 18 11 
150 310 30 200 9
-7 79 960 623
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
-7 79 960 623
9961490 0
0
6 Title:
5 Name:
0
0
0
13
11 Signal Gen~
195 240 443 0 19 64
0 0 0 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 1065353216
20
1 1000 0 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 832 0
5 -1/1V
-18 -30 17 -22
2 V1
-7 -40 7 -32
0
0
36 %D %1 %2 DC 0 SIN(0 1 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
8953 0 0
0
0
7 Ground~
168 274 461 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4441 0 0
0
0
7 Ground~
168 335 379 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3618 0 0
0
0
2 +V
167 439 447 0 1 3
0 4
0
0 0 54112 692
4 -15V
-4 -1 24 7
3 VEE
-1 7 20 15
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6153 0 0
0
0
2 +V
167 439 396 0 1 3
0 3
0
0 0 54112 0
3 15V
-11 -16 10 -8
3 VCC
-10 -27 11 -19
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5394 0 0
0
0
7 Ground~
168 385 479 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7734 0 0
0
0
10 Op-Amp5:A~
219 439 419 0 5 11
0 8 6 4 3 7
0
0 0 832 692
5 UA741
11 5 46 13
2 U3
13 -10 27 -2
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 256 1 0 0 0
1 U
9914 0 0
0
0
10 Capacitor~
219 329 452 0 2 5
0 7 5
0
0 0 832 90
5 1.6nF
11 -3 46 5
1 C
19 -12 26 -4
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3747 0 0
0
0
10 Capacitor~
219 385 452 0 2 5
0 2 8
0
0 0 832 90
5 1.6nF
10 -3 45 5
2 C1
14 -12 28 -4
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3549 0 0
0
0
9 Resistor~
219 354 425 0 2 5
0 5 8
0
0 0 864 0
3 10k
-10 -14 11 -6
1 R
-4 -24 3 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7931 0 0
0
0
9 Resistor~
219 445 357 0 2 5
0 6 7
0
0 0 864 0
6 3.694k
-22 -14 20 -6
2 R2
-8 -24 6 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9325 0 0
0
0
9 Resistor~
219 359 357 0 3 5
0 2 6 -1
0
0 0 864 0
6 6.306k
-21 -13 21 -5
2 R1
-8 -24 6 -16
6 3.694k
-21 -34 21 -26
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8903 0 0
0
0
9 Resistor~
219 300 424 0 3 5
0 2 5 -1
0
0 0 864 0
3 10k
-10 -14 11 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3834 0 0
0
0
14
2 1 0 0 0 0 0 1 2 0 0 3
271 448
274 448
274 455
1 1 0 0 0 0 0 1 13 0 0 4
271 438
274 438
274 424
282 424
1 4 3 0 0 4224 0 5 7 0 0 2
439 405
439 406
1 3 4 0 0 0 0 4 7 0 0 2
439 432
439 432
0 1 5 0 0 8192 0 0 10 14 0 3
328 424
328 425
336 425
2 0 6 0 0 8320 0 7 0 0 8 3
421 413
395 413
395 357
1 1 2 0 0 0 0 3 12 0 0 3
335 373
335 357
341 357
2 1 6 0 0 0 0 12 11 0 0 2
377 357
427 357
0 2 7 0 0 4096 0 0 11 10 0 3
490 419
490 357
463 357
1 5 7 0 0 8320 0 8 7 0 0 5
329 461
329 496
490 496
490 419
457 419
1 1 2 0 0 0 0 6 9 0 0 4
385 473
385 460
385 460
385 461
0 1 8 0 0 4224 0 0 7 13 0 2
385 425
421 425
2 2 8 0 0 0 0 10 9 0 0 3
372 425
385 425
385 443
2 2 5 0 0 8320 0 13 8 0 0 3
318 424
329 424
329 443
0
0
17 0 0
0
0
0
0 0 0
0
0 0 0
10 1 0.001 1e+009
0 0.0004 2e-006 2e-006
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
5049180 8550976 100 100 0 0
77 66 1217 606
170 222 1438 931
228 66
527 66
1217 66
1217 337
0 0
4.67281e-315 4.73699e-315 1.55453e-314 1.55453e-314 4.79266e-315 4.79266e-315
12441 0
4 0.0001 10
1
490 419
20 7 0 0 1	0 9 0 0
2688978 1341504 100 100 0 0
77 66 929 426
0 71 161 141
929 66
77 66
929 66
929 426
0 0
6.50121e-315 4.85009e-315 5.5705e-315 1.61805e-314 6.50121e-315 5.61194e-315
12385 0
4 5 10
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
