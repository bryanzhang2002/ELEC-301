CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 20 20 
10 13 13 10 20 13 20 20 14 20 
18 17 20 16 16 20 20 20 10 13 
20 18 11 
80 550 30 230 9
0 71 1920 515
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1920 515
9961490 256
0
6 Title:
5 Name:
0
0
0
17
7 Ground~
168 872 814 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8953 0 0
0
0
11 Signal Gen~
195 679 771 0 64 64
0 3 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 1065353216
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 1410949994
20
1 1000 0 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
5 -1/1V
-18 -30 17 -22
2 V2
-7 -40 7 -32
0
0
36 %D %1 %2 DC 0 SIN(0 1 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
4441 0 0
0
0
6 sxfer~
219 751 762 0 2 5
0 3 6
0
0 0 848 0
5 SXFER
-11 -31 24 -23
2 U1
0 -41 14 -33
0
0
11 %D %1 %2 %M
0
10 type:sxfer
0
5

0 0 0 0 0 0
65 0 0 0 1 0 0 0
1 U
3618 0 0
0
0
6 sxfer~
219 823 762 0 2 5
0 6 5
0
0 0 848 0
6 SXFER2
-14 -31 28 -23
2 U2
0 -41 14 -33
0
0
11 %D %1 %2 %M
0
10 type:sxfer
0
5

0 0 0 0 0 0
65 0 0 0 1 0 0 0
1 U
6153 0 0
0
0
6 sxfer~
219 895 762 0 2 5
0 5 4
0
0 0 848 0
6 SXFER3
-14 -31 28 -23
2 U3
0 -41 14 -33
0
0
11 %D %1 %2 %M
0
10 type:sxfer
0
5

0 0 0 0 0 0
65 0 0 0 1 0 0 0
1 U
5394 0 0
0
0
7 Ground~
168 409 708 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7734 0 0
0
0
10 Capacitor~
219 508 663 0 2 5
0 2 7
0
0 0 848 90
4 80pF
-38 0 -10 8
2 C3
-19 -10 -5 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
9914 0 0
0
0
10 Capacitor~
219 391 663 0 2 5
0 2 8
0
0 0 848 90
5 0.8nF
-40 6 -5 14
2 C2
-21 -11 -7 -3
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3747 0 0
0
0
10 Capacitor~
219 292 663 0 2 5
0 2 9
0
0 0 848 90
3 8nF
-26 3 -5 11
2 C1
-23 -8 -9 0
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3549 0 0
0
0
11 Signal Gen~
195 193 663 0 64 64
0 10 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 1065353216
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 -1258556724
20
1 1000 0 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
5 -1/1V
-18 -30 17 -22
2 V1
-7 -40 7 -32
0
0
36 %D %1 %2 DC 0 SIN(0 1 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
7931 0 0
0
0
9 Resistor~
219 944 787 0 3 5
0 2 4 -1
0
0 0 880 90
3 500
5 0 26 8
2 R6
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9325 0 0
0
0
9 Resistor~
219 526 663 0 3 5
0 2 7 -1
0
0 0 880 90
3 500
6 0 27 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8903 0 0
0
0
9 Resistor~
219 409 663 0 3 5
0 2 8 -1
0
0 0 880 90
2 1k
8 0 22 8
2 R5
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3834 0 0
0
0
9 Resistor~
219 310 663 0 3 5
0 2 9 -1
0
0 0 880 90
2 1k
8 0 22 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3363 0 0
0
0
9 Resistor~
219 454 636 0 2 5
0 8 7
0
0 0 880 0
3 500
-10 -14 11 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7668 0 0
0
0
9 Resistor~
219 355 636 0 2 5
0 9 8
0
0 0 880 0
3 500
-10 -14 11 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4718 0 0
0
0
9 Resistor~
219 247 636 0 2 5
0 10 9
0
0 0 880 0
3 500
-10 -13 11 -5
2 R7
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3874 0 0
0
0
22
1 1 3 0 0 8320 0 2 3 0 0 3
710 766
710 762
727 762
1 2 2 0 0 8192 0 1 2 0 0 4
872 808
872 806
710 806
710 776
1 1 2 0 0 0 0 11 1 0 0 4
944 805
944 806
872 806
872 808
2 2 4 0 0 4224 0 5 11 0 0 3
933 762
944 762
944 769
2 1 5 0 0 4224 0 4 5 0 0 4
861 762
876 762
876 762
871 762
2 1 6 0 0 4224 0 3 4 0 0 4
789 762
813 762
813 762
799 762
1 0 2 0 0 0 0 6 0 0 12 2
409 702
409 691
1 0 2 0 0 0 0 7 0 0 13 2
508 672
508 691
1 0 2 0 0 0 0 14 0 0 13 2
310 681
310 691
2 0 2 0 0 0 0 10 0 0 13 4
224 668
226 668
226 691
292 691
1 0 2 0 0 0 0 8 0 0 13 2
391 672
391 691
1 0 2 0 0 0 0 13 0 0 13 2
409 681
409 691
1 1 2 0 0 8320 0 9 12 0 0 4
292 672
292 691
526 691
526 681
2 0 7 0 0 4096 0 7 0 0 15 2
508 654
508 636
2 2 7 0 0 4224 0 15 12 0 0 3
472 636
526 636
526 645
2 0 8 0 0 4096 0 13 0 0 18 2
409 645
409 636
2 0 8 0 0 4096 0 8 0 0 18 2
391 654
391 636
2 1 8 0 0 4224 0 16 15 0 0 2
373 636
436 636
2 0 9 0 0 4096 0 14 0 0 21 2
310 645
310 637
2 0 9 0 0 4096 0 9 0 0 21 2
292 654
292 637
2 1 9 0 0 8320 0 17 16 0 0 4
265 636
265 637
337 637
337 636
1 1 10 0 0 4224 0 10 17 0 0 3
224 658
224 636
229 636
0
0
8 0 0
0
0
0
0 0 0
0
0 0 0
10 1 1 1e+009
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
460566 4290624 100 100 0 0
77 66 1886 426
-74 492 1846 1013
1886 66
77 66
1886 66
1886 336
0 0
1e+009 1 0 -180 1e+009 1e+009
12435 0
4 3e+008 5e+008
1
514 636
0 7 0 0 1	0 15 0 0
3082998 8419904 100 100 0 0
77 66 917 396
960 71 1920 551
917 66
77 66
917 66
917 396
0 0
0 0 0 0 0 0
12409 0
4 0.001 0.5
0
4524378 272791618 100 100 0 0
77 66 1889 396
0 551 1920 1031
1886 66
77 66
1889 87
1889 182
0 0
0 0 0 0 0 0
45299 0
4 300000 500000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
