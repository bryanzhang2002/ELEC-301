CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 20 20 
10 13 13 10 20 13 20 20 14 20 
18 17 20 16 16 20 20 20 10 13 
20 18 11 
620 180 30 200 9
82 122 1906 1013
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
82 122 1906 1013
77070354 256
0
6 Title:
5 Name:
0
0
0
7
12 NPN Trans:B~
219 738 423 0 3 7
0 3 5 4
0
0 0 848 0
6 2N4401
18 0 60 8
2 Q1
32 -10 46 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
8953 0 0
0
0
7 Ground~
168 729 495 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4441 0 0
0
0
2 +V
167 729 342 0 1 3
0 6
0
0 0 54128 0
3 15V
-9 -15 12 -7
3 VCC
-9 -25 12 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3618 0 0
0
0
9 Resistor~
219 747 468 0 3 5
0 2 4 -1
0
0 0 880 90
4 4.3k
15 6 43 14
2 RE
7 -5 21 3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6153 0 0
0
0
9 Resistor~
219 702 468 0 3 5
0 2 5 -1
0
0 0 880 90
3 62k
-39 5 -18 13
3 RB2
-30 -8 -9 0
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5394 0 0
0
0
9 Resistor~
219 702 378 0 4 5
0 5 6 0 1
0
0 0 880 90
4 110k
-41 6 -13 14
3 RB1
-27 -5 -6 3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7734 0 0
0
0
9 Resistor~
219 747 378 0 4 5
0 3 6 0 1
0
0 0 880 90
4 5.1k
5 6 33 14
2 RC
8 -5 22 3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9914 0 0
0
0
8
1 1 3 0 0 4224 0 1 7 0 0 3
743 405
743 396
747 396
3 2 4 0 0 4224 0 1 4 0 0 3
743 441
743 450
747 450
1 1 2 0 0 4096 0 2 4 0 0 3
729 489
747 489
747 486
1 1 2 0 0 8320 0 5 2 0 0 3
702 486
702 489
729 489
0 2 5 0 0 4224 0 0 5 6 0 2
702 423
702 450
1 2 5 0 0 0 0 6 1 0 0 3
702 396
702 423
720 423
1 2 6 0 0 4224 0 3 6 0 0 3
729 351
702 351
702 360
2 1 6 0 0 0 0 7 3 0 0 3
747 360
747 351
729 351
0
0
1 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
723446 1079360 100 100 0 0
0 0 0 0
39 102 200 172
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12401 0
4 3 10
1
743 446
0 4 0 0 1	0 2 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
