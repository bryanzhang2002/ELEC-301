CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 20 20 
10 13 13 10 20 13 20 20 14 20 
18 17 20 16 16 20 20 20 10 13 
20 18 11 
330 270 30 200 9
0 71 1440 791
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1440 791
77070354 256
0
6 Title:
5 Name:
0
0
0
11
7 Ground~
168 720 477 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8953 0 0
0
0
10 Capacitor~
219 837 396 0 2 5
0 3 5
0
0 0 848 0
3 1uF
-11 -18 10 -10
2 C4
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
4441 0 0
0
0
10 Capacitor~
219 702 396 0 2 5
0 4 3
0
0 0 848 0
3 2pF
-11 -18 10 -10
2 C3
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3618 0 0
0
0
12 V->I Source~
200 702 432 0 4 9
0 3 2 4 2
0
0 0 17232 0
3 0.1
46 1 67 9
5 VcIs1
39 -9 74 -1
0
0
17 %D %1 %2 %3 %4 %V
0
0
0
9

0 3 4 1 2 3 4 1 2 0
71 0 0 0 0 0 0 0
4 VcIs
6153 0 0
0
0
10 Capacitor~
219 621 423 0 2 5
0 2 4
0
0 0 848 90
4 10pF
8 0 36 8
2 C2
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5394 0 0
0
0
10 Capacitor~
219 567 396 0 2 5
0 6 4
0
0 0 848 0
3 1uF
-11 -18 10 -10
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7734 0 0
0
0
11 Signal Gen~
195 468 423 0 19 64
0 7 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 1065353216
20
1 1000 0 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
5 -1/1V
-18 -30 17 -22
2 V1
-7 -40 7 -32
0
0
36 %D %1 %2 DC 0 SIN(0 1 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
9914 0 0
0
0
9 Resistor~
219 873 423 0 3 5
0 2 5 -1
0
0 0 880 90
2 4k
8 0 22 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3747 0 0
0
0
9 Resistor~
219 801 423 0 3 5
0 2 3 -1
0
0 0 880 90
2 4k
8 0 22 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3549 0 0
0
0
9 Resistor~
219 585 423 0 3 5
0 2 4 -1
0
0 0 880 90
2 1k
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7931 0 0
0
0
9 Resistor~
219 531 396 0 2 5
0 7 6
0
0 0 880 0
2 50
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9325 0 0
0
0
17
4 0 2 0 0 4096 0 4 0 0 9 2
682 459
682 471
2 1 2 0 0 0 0 4 1 0 0 3
722 459
720 459
720 471
1 0 2 0 0 4096 0 9 0 0 4 2
801 441
801 471
1 1 2 0 0 4096 0 1 8 0 0 3
720 471
873 471
873 441
1 0 3 0 0 4096 0 4 0 0 12 2
722 405
722 396
3 0 4 0 0 4096 0 4 0 0 15 2
682 405
682 396
1 0 2 0 0 0 0 5 0 0 9 2
621 432
621 471
1 0 2 0 0 0 0 10 0 0 9 2
585 441
585 471
2 1 2 0 0 12416 0 7 1 0 0 4
499 428
504 428
504 471
720 471
2 2 5 0 0 4224 0 2 8 0 0 3
846 396
873 396
873 405
2 0 3 0 0 0 0 9 0 0 12 2
801 405
801 396
2 1 3 0 0 4224 0 3 2 0 0 2
711 396
828 396
2 0 4 0 0 0 0 10 0 0 15 2
585 405
585 396
2 0 4 0 0 4096 0 5 0 0 15 2
621 414
621 396
2 1 4 0 0 4224 0 6 3 0 0 2
576 396
693 396
2 1 6 0 0 4224 0 11 6 0 0 2
549 396
558 396
1 1 7 0 0 8320 0 7 11 0 0 4
499 418
504 418
504 396
513 396
0
0
8 0 0
0
0
0
0 0 0
0
0 0 0
10 1 0.01 1e+011
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
1836116 4290624 100 100 0 0
77 66 1884 876
0 71 1920 1032
1300 66
661 66
1884 130
1884 144
0 0
6.2887e+006 159.015 45.7778 42.7875 1e+011 1e+011
12307 0
5 3e+010 5e+010
1
867 396
20 5 0 0 1	0 10 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
