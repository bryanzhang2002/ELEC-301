CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 20 20 
10 13 13 10 20 13 20 20 14 20 
18 17 20 16 16 20 20 20 10 13 
20 18 11 
380 220 30 200 9
-595 259 1325 1072
7 5.000 V
7 5.000 V
3 GND
0 0
24 133.333 0 1 1
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
-595 259 1325 1072
76546066 256
0
6 Title:
5 Name:
0
0
0
4
7 Ground~
168 819 378 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8953 0 0
0
0
9 V Source~
197 900 351 0 2 5
0 3 2
0
0 0 17264 0
2 5V
16 0 30 8
3 Vce
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
4441 0 0
0
0
9 V Source~
197 747 351 0 2 5
0 4 2
0
0 0 17008 0
3 10V
13 0 34 8
3 Vbe
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
3618 0 0
0
0
12 NPN Trans:B~
219 810 324 0 3 7
0 3 4 2
0
0 0 848 0
6 2N3904
18 0 60 8
2 Q1
32 -10 46 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
6153 0 0
0
0
5
1 0 2 0 0 0 0 1 0 0 5 2
819 372
819 372
1 1 3 0 0 4224 0 4 2 0 0 3
815 306
900 306
900 330
1 2 4 0 0 8320 0 3 4 0 0 3
747 330
747 324
792 324
3 0 2 0 0 4112 0 4 0 0 5 2
815 342
815 372
2 2 2 0 0 4224 0 3 2 0 0 2
747 372
900 372
0
0
5 0 0
0
0
3 Vbe
0 0.7 0.01
0
0 0 0
3 0 1 4
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
592290 1210432 100 100 0 0
0 0 0 0
0 71 161 141
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 2 5e+035
0
592278 2255424 100 100 0 0
77 66 977 336
814 316 1825 733
976 66
77 66
977 66
977 336
0 0
0.7 0 4.5e-005 -9e-006 0.7 0.7
12441 0
4 0.2 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
