CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 20 20 
10 13 13 10 20 13 20 20 14 20 
18 17 20 16 16 20 20 20 10 13 
20 18 11 
0 190 30 260 9
0 71 1920 915
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1920 915
9961490 0
0
6 Title:
5 Name:
0
0
0
17
7 Ground~
168 174 367 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8953 0 0
0
0
7 Ground~
168 282 450 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4441 0 0
0
0
7 Ground~
168 184 448 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3618 0 0
0
0
10 Capacitor~
219 250 393 0 2 5
0 9 10
0
0 0 848 0
4 10uF
-14 -18 14 -10
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6153 0 0
0
0
2 +V
167 333 425 0 1 3
0 11
0
0 0 54128 180
3 -5V
6 -2 27 6
3 VEE
7 -12 28 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
5394 0 0
0
0
12 NPN Trans:B~
219 328 393 0 3 7
0 12 10 11
0
0 0 848 0
6 2N3904
18 0 60 8
2 Q3
32 -10 46 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
7734 0 0
0
0
7 Ground~
168 410 326 0 1 3
0 2
0
0 0 53360 90
0
4 GND1
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9914 0 0
0
0
12 NPN Trans:B~
219 391 327 0 3 7
0 3 2 12
0
0 0 848 512
6 2N3904
-64 0 -22 8
2 Q2
-50 -10 -36 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
3747 0 0
0
0
12 NPN Trans:B~
219 265 327 0 3 7
0 5 6 12
0
0 0 848 0
6 2N3904
18 0 60 8
2 Q1
32 -10 46 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
3549 0 0
0
0
2 +V
167 326 224 0 1 3
0 4
0
0 0 54128 0
2 5V
-6 -12 8 -4
3 Vcc
-10 -22 11 -14
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
7931 0 0
0
0
11 Signal Gen~
195 143 426 0 24 64
0 8 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1148846079 -1115349319 1032134329
0 814313567 814313567 973279855 981668463
20
0 1000 -0.065 0.065 0 1e-009 1e-009 0.0005 0.001 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
9 -65m/65mV
-32 -30 31 -22
2 V2
-7 -40 7 -32
0
0
45 %D %1 %2 DC 0 PULSE(-65m 65m 0 1n 1n 500u 1m)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
9325 0 0
0
0
11 Signal Gen~
195 139 340 0 19 64
0 7 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1203982336 0 1028443341
20
1 100000 0 0.05 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
9 -50m/50mV
-32 -30 31 -22
2 V1
-7 -40 7 -32
0
0
40 %D %1 %2 DC 0 SIN(0 50m 100k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
8903 0 0
0
0
9 Resistor~
219 206 393 0 2 5
0 8 9
0
0 0 880 0
2 2k
-7 -14 7 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3834 0 0
0
0
9 Resistor~
219 282 423 0 3 5
0 2 10 -1
0
0 0 880 90
4 200k
3 0 31 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3363 0 0
0
0
9 Resistor~
219 381 270 0 4 5
0 3 4 0 1
0
0 0 880 90
2 1k
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7668 0 0
0
0
9 Resistor~
219 270 268 0 4 5
0 5 4 0 1
0
0 0 880 90
2 1k
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4718 0 0
0
0
9 Resistor~
219 212 327 0 2 5
0 7 6
0
0 0 880 0
2 50
-7 -14 7 -6
2 Rs
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3874 0 0
0
0
17
1 2 2 0 0 4224 0 1 12 0 0 3
174 361
174 345
170 345
1 1 2 0 0 0 0 2 14 0 0 4
282 444
282 440
282 440
282 441
1 1 3 0 0 8320 0 8 15 0 0 3
382 309
381 309
381 288
1 2 4 0 0 8192 0 10 15 0 0 4
326 233
326 241
381 241
381 252
2 1 4 0 0 8320 0 16 10 0 0 4
270 250
270 241
326 241
326 233
1 1 5 0 0 4224 0 9 16 0 0 2
270 309
270 286
2 2 6 0 0 4224 0 17 9 0 0 2
230 327
247 327
1 1 7 0 0 12416 0 12 17 0 0 4
170 335
174 335
174 327
194 327
2 1 2 0 0 128 0 11 3 0 0 3
174 431
184 431
184 442
1 1 8 0 0 8320 0 11 13 0 0 4
174 421
180 421
180 393
188 393
2 1 9 0 0 4224 0 13 4 0 0 2
224 393
241 393
0 2 10 0 0 4096 0 0 14 13 0 2
282 393
282 405
2 2 10 0 0 4224 0 4 6 0 0 2
259 393
310 393
1 3 11 0 0 4224 0 5 6 0 0 2
333 410
333 411
1 0 12 0 0 4096 0 6 0 0 16 2
333 375
333 353
3 3 12 0 0 8320 0 9 8 0 0 4
270 345
270 353
382 353
382 345
1 2 2 0 0 0 0 7 8 0 0 4
403 327
409 327
409 327
405 327
0
0
16 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 1e-006 1e-006
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
6556592 8419904 100 100 0 0
77 66 1877 876
0 71 1920 1032
1874 66
77 66
1877 66
1877 876
381 300
0.00499167 0 8 -4 0.005 0.005
12297 0
4 0.001 3
1
270 303
20 5 0 0 1	0 6 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
