CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 20 20 
10 13 13 10 20 13 20 20 14 20 
18 17 20 16 16 20 20 20 10 13 
20 18 11 
170 250 30 400 9
0 71 1920 1028
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1920 1028
77070354 256
0
6 Title:
5 Name:
0
0
0
8
10 Capacitor~
219 513 351 0 1 5
0 0
0
0 0 576 0
3 1uF
-11 -18 10 -10
2 C3
-7 -21 7 -13
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
8953 0 0
0
0
7 Ground~
168 441 387 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 512 0 0 0 0
3 GND
4441 0 0
0
0
7 Ground~
168 396 387 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3618 0 0
0
0
7 Ground~
168 540 387 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
6153 0 0
0
0
9 Resistor~
219 540 369 0 3 5
0 2 3 -1
0
0 0 864 90
2 1k
8 0 22 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5394 0 0
0
0
9 Resistor~
219 468 351 0 2 5
0 4 3
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7734 0 0
0
0
9 Resistor~
219 441 369 0 2 5
0 6 4
0
0 0 880 90
2 1k
8 1 22 9
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 512 1 0 0 0
1 R
9914 0 0
0
0
9 Resistor~
219 414 351 0 3 5
0 2 5 -1
0
0 0 880 0
2 50
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3747 0 0
0
0
7
2 2 0 0 0 0 0 1 5 0 0 2
522 351
540 351
2 1 0 0 0 0 0 6 1 0 0 2
486 351
504 351
2 2 0 0 0 0 0 8 7 0 0 2
432 351
441 351
1 2 0 0 0 0 0 6 7 0 0 2
450 351
441 351
1 1 0 0 0 0 0 2 7 0 0 2
441 381
441 387
1 1 2 0 0 4096 0 4 5 0 0 2
540 381
540 387
1 1 2 0 0 8320 0 8 3 0 0 2
396 351
396 381
0
0
8 0 0
0
0
0
0 0 0
0
0 0 0
10 1 0.01 1e+009
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
1444030 4290624 100 100 0 0
77 66 1881 876
0 71 1920 1032
1881 66
601 66
1881 231
1881 244
0 0
1e+009 15.6719 -6.66667 -9.55556 1e+009 1e+009
12435 2
5 3e+008 5e+008
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
