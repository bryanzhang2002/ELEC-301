CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 20 20 
10 13 13 10 20 13 20 20 14 20 
18 17 20 16 16 20 20 20 10 13 
20 18 11 
90 390 30 400 9
48 106 1872 997
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
48 106 1872 997
76021778 256
0
6 Title:
5 Name:
0
0
0
18
7 Ground~
168 126 459 0 1 3
0 0
0
0 0 53344 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8953 0 0
0
0
7 Ground~
168 504 450 0 1 3
0 0
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4441 0 0
0
0
7 Ground~
168 441 450 0 1 3
0 0
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3618 0 0
0
0
7 Ground~
168 198 450 0 1 3
0 0
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
6153 0 0
0
0
9 Resistor~
219 504 423 0 1 5
0 0
0
0 0 864 90
4 5.1k
4 2 32 10
2 RL
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5394 0 0
0
0
10 Capacitor~
219 477 405 0 1 5
0 0
0
0 0 832 0
4 10uF
-14 -18 14 -10
3 CC2
-10 -28 11 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7734 0 0
0
0
9 Resistor~
219 441 423 0 1 5
0 0
0
0 0 864 90
4 5.1k
5 2 33 10
2 RC
6 -8 20 0
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9914 0 0
0
0
7 Ground~
168 297 522 0 1 3
0 0
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3747 0 0
0
0
10 Capacitor~
219 315 495 0 1 5
0 0
0
0 0 832 90
4 10uF
8 0 36 8
2 CE
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3549 0 0
0
0
9 Resistor~
219 279 495 0 1 5
0 0
0
0 0 864 90
4 4.3k
-33 1 -5 9
2 RE
-20 -10 -6 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7931 0 0
0
0
12 V->I Source~
200 378 432 0 1 9
0 0
0
0 0 16704 0
4 0.04
-12 -17 16 -9
5 gmvpi
39 -9 74 -1
0
0
17 %D %1 %2 %3 %4 %V
0
0
0
9

0 3 4 1 2 3 4 1 2 0
71 0 0 0 0 0 0 0
4 VcIs
9325 0 0
0
0
10 Capacitor~
219 378 396 0 1 5
0 0
0
0 0 832 0
3 1uF
-11 -18 10 -10
2 Cu
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
8903 0 0
0
0
10 Capacitor~
219 297 432 0 1 5
0 0
0
0 0 832 90
4 25pF
9 2 37 10
3 Cpi
8 -11 29 -3
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3834 0 0
0
0
9 Resistor~
219 243 432 0 1 5
0 0
0
0 0 864 90
5 2.95k
4 1 39 9
3 Rpi
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3363 0 0
0
0
9 Resistor~
219 198 432 0 1 5
0 0
0
0 0 864 90
5 39.7k
3 0 38 8
3 RBB
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7668 0 0
0
0
10 Capacitor~
219 180 405 0 1 5
0 0
0
0 0 832 0
4 10uF
-14 -18 14 -10
3 CC1
-10 -28 11 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
4718 0 0
0
0
9 Resistor~
219 144 405 0 1 5
0 0
0
0 0 864 0
2 50
-7 -14 7 -6
2 Rs
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3874 0 0
0
0
11 Signal Gen~
195 90 441 0 19 64
0 0 0 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 1065353216
20
1 1000 0 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 832 0
5 -1/1V
-18 -30 17 -22
2 V1
-7 -40 7 -32
0
0
36 %D %1 %2 DC 0 SIN(0 1 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
6671 0 0
0
0
20
2 0 0 0 0 0 0 13 0 0 17 2
297 423
297 405
2 0 0 0 0 0 0 15 0 0 18 2
198 414
198 405
2 4 0 0 0 0 0 11 11 0 0 2
398 459
358 459
2 1 0 0 0 0 0 18 1 0 0 3
121 446
126 446
126 453
1 1 0 0 0 0 0 2 5 0 0 4
504 444
504 447
504 447
504 441
1 1 0 0 0 0 0 3 7 0 0 4
441 444
441 447
441 447
441 441
2 2 0 0 0 0 0 6 5 0 0 2
486 405
504 405
1 1 0 0 0 0 0 11 6 0 0 2
398 405
468 405
1 1 0 0 0 0 0 9 8 0 0 3
315 504
315 516
297 516
1 1 0 0 0 0 0 10 8 0 0 3
279 513
279 516
297 516
0 2 0 0 0 0 0 0 9 12 0 3
297 477
315 477
315 486
1 2 0 0 0 16 0 13 10 0 0 3
297 441
297 477
279 477
1 4 0 0 0 0 0 14 11 0 0 3
243 450
243 459
358 459
1 1 0 0 0 0 0 4 15 0 0 2
198 444
198 450
2 1 0 0 0 0 0 12 11 0 0 3
387 396
398 396
398 405
1 3 0 0 0 0 0 12 11 0 0 3
369 396
358 396
358 405
0 3 0 0 0 0 0 0 11 18 0 2
243 405
358 405
2 2 0 0 0 0 0 16 14 0 0 3
189 405
243 405
243 414
2 1 0 0 0 0 0 17 16 0 0 4
162 405
177 405
177 405
171 405
1 1 0 0 0 0 0 18 17 0 0 3
121 436
121 405
126 405
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 100 100 0 0
77 66 1001 516
0 0 0 0
1001 66
77 66
1001 66
1001 516
0 0
1e+011 0.001 80 -160 1e+011 1e+011
12435 4
0 30 50
0
0 0 100 100 0 0
77 66 1889 396
0 0 0 0
1889 66
77 66
1889 66
1889 396
0 0
100 1 18 0 99 99
12307 0
0 30 50
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
